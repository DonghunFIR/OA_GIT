----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 2024/01/31 11:39:21
-- Design Name: 
-- Module Name: Digital_Potentiometer - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Digital_Potentiometer is
	Port ( 
	--===== INPUT =====--
	-- CLOCK --
	m_sys_clk_160M			: in std_logic;
	
	);
end Digital_Potentiometer;

architecture Behavioral of Digital_Potentiometer is
--
---
begin
---
--

end Behavioral;
